// example Verilog code with AND Gate
module and_verrilog(a, b, c);
   input a, b;
   output c;
   assign c = a & b;
endmodule